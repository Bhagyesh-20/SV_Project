interface intf;
  
  logic [3:0] A_mag;
  logic [3:0] B_mag;
  logic       A_sign;
  logic       B_sign;
  logic [4:0] Out_mag;     
  logic       Out_sign;  

endinterface
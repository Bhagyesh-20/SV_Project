interface intf;
  
  logic [7:0] a;
  logic [7:0] b; 
  logic sign_a; 
  logic sign_b;
  logic  sign;
  logic  [8:0] result;
  
endinterface
class enviroment;
endclass